// *!***************************************************************************
// *! Copyright 2019 International Business Machines
// *!
// *! Licensed under the Apache License, Version 2.0 (the "License");
// *! you may not use this file except in compliance with the License.
// *! You may obtain a copy of the License at
// *! http://www.apache.org/licenses/LICENSE-2.0 
// *!
// *! The patent license granted to you in Section 3 of the License, as applied
// *! to the "Work," hereby includes implementations of the Work in physical form. 
// *!
// *! Unless required by applicable law or agreed to in writing, the reference design
// *! distributed under the License is distributed on an "AS IS" BASIS,
// *! WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// *! See the License for the specific language governing permissions and
// *! limitations under the License.
// *!***************************************************************************
module base_ademux#
  (
   parameter ways = 2
   )
  (
   input [0:ways-1]   sel,
   input 	      i_v,
   output 	      i_r,
   output [0:ways-1]  o_v,
   input [0:ways-1]   o_r
   );

   assign i_r = &(~sel | o_r);
   assign o_v = sel & {ways{i_v}};
endmodule // base_mux
   
		
