// *!***************************************************************************
// *! Copyright 2019 International Business Machines
// *!
// *! Licensed under the Apache License, Version 2.0 (the "License");
// *! you may not use this file except in compliance with the License.
// *! You may obtain a copy of the License at
// *! http://www.apache.org/licenses/LICENSE-2.0 
// *!
// *! The patent license granted to you in Section 3 of the License, as applied
// *! to the "Work," hereby includes implementations of the Work in physical form. 
// *!
// *! Unless required by applicable law or agreed to in writing, the reference design
// *! distributed under the License is distributed on an "AS IS" BASIS,
// *! WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// *! See the License for the specific language governing permissions and
// *! limitations under the License.
// *!***************************************************************************
module base_vlat (clk, reset, din, q);
   parameter width=1;
   parameter [width-1:0] rstv = 0;
   input clk;
   input reset;
   input [width-1:0] din;
   output [width-1:0] q;
   reg [width-1:0]    q_int;

   initial q_int = rstv;

   always@(posedge clk or posedge reset)
     if (reset) q_int <= rstv;
     else q_int <= din;
   assign q = q_int;
   
endmodule // base_vlat


   
  
