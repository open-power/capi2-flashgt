// *!***************************************************************************
// *! Copyright 2019 International Business Machines
// *!
// *! Licensed under the Apache License, Version 2.0 (the "License");
// *! you may not use this file except in compliance with the License.
// *! You may obtain a copy of the License at
// *! http://www.apache.org/licenses/LICENSE-2.0 
// *!
// *! The patent license granted to you in Section 3 of the License, as applied
// *! to the "Work," hereby includes implementations of the Work in physical form. 
// *!
// *! Unless required by applicable law or agreed to in writing, the reference design
// *! distributed under the License is distributed on an "AS IS" BASIS,
// *! WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// *! See the License for the specific language governing permissions and
// *! limitations under the License.
// *!***************************************************************************
module ktms_afu_errmux#(parameter rc_width=1)
   (input i_ok,
    input [0:rc_width-1] i_rc,
    input i_err,
    input [0:rc_width-1] i_err_rc,
    output o_ok,
    output [0:rc_width-1] o_rc
    );
   assign o_ok = i_ok & ~i_err;
   assign o_rc = i_ok ? (i_err ? i_err_rc : {rc_width{1'b0}}) : i_rc;
endmodule // ktms_afu_errmux

