// *!***************************************************************************
// *! Copyright 2019 International Business Machines
// *!
// *! Licensed under the Apache License, Version 2.0 (the "License");
// *! you may not use this file except in compliance with the License.
// *! You may obtain a copy of the License at
// *! http://www.apache.org/licenses/LICENSE-2.0 
// *!
// *! The patent license granted to you in Section 3 of the License, as applied
// *! to the "Work," hereby includes implementations of the Work in physical form. 
// *!
// *! Unless required by applicable law or agreed to in writing, the reference design
// *! distributed under the License is distributed on an "AS IS" BASIS,
// *! WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// *! See the License for the specific language governing permissions and
// *! limitations under the License.
// *!***************************************************************************
module capi_parity_gen#(parameter dwidth=64, parameter width=2)
   (input [0:dwidth*width-1] i_d,
    output [0:width-1] o_d
    );

   genvar 	       i;
   generate
      for(i=0; i<width; i=i+1)
	begin :gen
	   assign o_d[i] = ~(^(i_d[i*dwidth:((i+1)*dwidth)-1]));
	end
   endgenerate
endmodule // capi_parity_gen

   
  
    
					    
